library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity winner_rom is
   Port (
       x_coord : in std_logic_vector(6 downto 0);
	   y_coord : in std_logic_vector(5 downto 0);
       rgb : out std_logic_vector(5 downto 0)
   );
end winner_rom;


architecture Behavioral of winner_rom is
signal total : std_logic_vector(12 downto 0);

begin
total <= y_coord & x_coord;
   process(total)
   begin
	case total is
		when "0100111000010" => rgb <= "000000";
        when "0100111000011" => rgb <= "000000";
        when "0100111000100" => rgb <= "000000";
        when "0100111000101" => rgb <= "000000";
        when "0101000110111" => rgb <= "000000";
        when "0101000111000" => rgb <= "000000";
        when "0101000111001" => rgb <= "000000";
        when "0101000111010" => rgb <= "000000";
        when "0101000111011" => rgb <= "000000";
        when "0101000111100" => rgb <= "000000";
        when "0101000111101" => rgb <= "000000";
        when "0101001000000" => rgb <= "000000";
        when "0101001000001" => rgb <= "000000";
        when "0101001000010" => rgb <= "000000";
        when "0101001000011" => rgb <= "100000";
        when "0101001000100" => rgb <= "100000";
        when "0101001000101" => rgb <= "100000";
        when "0101001000110" => rgb <= "000000";
        when "0101001000111" => rgb <= "000000";
        when "0101001001011" => rgb <= "000000";
        when "0101001001100" => rgb <= "000000";
        when "0101001001101" => rgb <= "000000";
        when "0101010000010" => rgb <= "000000";
        when "0101010000011" => rgb <= "000000";
        when "0101010010010" => rgb <= "000000";
        when "0101010010011" => rgb <= "000000";
        when "0101010010100" => rgb <= "000000";
        when "0101010010101" => rgb <= "000000";
        when "0101010010110" => rgb <= "000000";
        when "0101010011010" => rgb <= "000000";
        when "0101010011011" => rgb <= "000000";
        when "0101010011100" => rgb <= "000000";
        when "0101010011101" => rgb <= "000000";
        when "0101010011110" => rgb <= "000000";
        when "0101010100100" => rgb <= "000000";
        when "0101010100101" => rgb <= "000000";
        when "0101010100110" => rgb <= "000000";
        when "0101010100111" => rgb <= "000000";
        when "0101010101000" => rgb <= "000000";
        when "0101010101001" => rgb <= "000000";
        when "0101010101010" => rgb <= "000000";
        when "0101010101011" => rgb <= "000000";
        when "0101010101100" => rgb <= "000000";
        when "0101010110010" => rgb <= "000000";
        when "0101010110011" => rgb <= "000000";
        when "0101010110100" => rgb <= "000000";
        when "0101010110101" => rgb <= "000000";
        when "0101010110110" => rgb <= "000000";
        when "0101010110111" => rgb <= "000000";
        when "0101010111000" => rgb <= "100110";
        when "0101010111001" => rgb <= "100110";
        when "0101010111010" => rgb <= "100110";
        when "0101010111011" => rgb <= "100110";
        when "0101010111100" => rgb <= "100110";
        when "0101010111101" => rgb <= "000000";
        when "0101010111110" => rgb <= "000000";
        when "0101010111111" => rgb <= "000000";
        when "0101011000000" => rgb <= "000000";
        when "0101011000001" => rgb <= "100000";
        when "0101011000010" => rgb <= "100000";
        when "0101011000011" => rgb <= "100000";
        when "0101011000100" => rgb <= "100000";
        when "0101011000101" => rgb <= "100000";
        when "0101011000110" => rgb <= "100000";
        when "0101011000111" => rgb <= "000000";
        when "0101011001000" => rgb <= "000000";
        when "0101011001010" => rgb <= "000000";
        when "0101011001011" => rgb <= "101000";
        when "0101011001100" => rgb <= "101000";
        when "0101011001101" => rgb <= "000000";
        when "0101100000001" => rgb <= "000000";
        when "0101100000010" => rgb <= "100000";
        when "0101100000011" => rgb <= "000000";
        when "0101100010001" => rgb <= "000000";
        when "0101100010010" => rgb <= "000000";
        when "0101100010011" => rgb <= "100000";
        when "0101100010100" => rgb <= "100000";
        when "0101100010101" => rgb <= "100000";
        when "0101100010110" => rgb <= "000000";
        when "0101100010111" => rgb <= "000000";
        when "0101100011000" => rgb <= "000000";
        when "0101100011001" => rgb <= "000000";
        when "0101100011010" => rgb <= "000000";
        when "0101100011011" => rgb <= "000000";
        when "0101100011100" => rgb <= "000000";
        when "0101100011101" => rgb <= "101000";
        when "0101100011110" => rgb <= "101000";
        when "0101100011111" => rgb <= "000000";
        when "0101100100100" => rgb <= "000000";
        when "0101100100101" => rgb <= "101000";
        when "0101100100110" => rgb <= "101000";
        when "0101100100111" => rgb <= "101000";
        when "0101100101000" => rgb <= "000000";
        when "0101100101001" => rgb <= "001010";
        when "0101100101010" => rgb <= "001010";
        when "0101100101011" => rgb <= "001010";
        when "0101100101100" => rgb <= "000000";
        when "0101100101101" => rgb <= "000000";
        when "0101100110010" => rgb <= "000000";
        when "0101100110011" => rgb <= "001010";
        when "0101100110100" => rgb <= "001010";
        when "0101100110101" => rgb <= "001010";
        when "0101100110110" => rgb <= "000000";
        when "0101100110111" => rgb <= "100110";
        when "0101100111000" => rgb <= "100110";
        when "0101100111001" => rgb <= "100110";
        when "0101100111010" => rgb <= "100110";
        when "0101100111011" => rgb <= "100110";
        when "0101100111100" => rgb <= "100110";
        when "0101100111101" => rgb <= "100110";
        when "0101100111110" => rgb <= "100110";
        when "0101100111111" => rgb <= "100110";
        when "0101101000000" => rgb <= "100110";
        when "0101101000001" => rgb <= "000000";
        when "0101101000010" => rgb <= "100000";
        when "0101101000011" => rgb <= "100000";
        when "0101101000100" => rgb <= "100000";
        when "0101101000101" => rgb <= "100000";
        when "0101101000110" => rgb <= "100000";
        when "0101101000111" => rgb <= "100000";
        when "0101101001000" => rgb <= "100000";
        when "0101101001001" => rgb <= "000000";
        when "0101101001010" => rgb <= "000000";
        when "0101101001011" => rgb <= "000000";
        when "0101101001100" => rgb <= "101000";
        when "0101101001101" => rgb <= "000000";
        when "0101110000001" => rgb <= "000000";
        when "0101110000010" => rgb <= "100000";
        when "0101110000011" => rgb <= "100000";
        when "0101110000100" => rgb <= "000000";
        when "0101110000101" => rgb <= "000000";
        when "0101110010001" => rgb <= "000000";
        when "0101110010010" => rgb <= "100000";
        when "0101110010011" => rgb <= "100000";
        when "0101110010100" => rgb <= "100000";
        when "0101110010101" => rgb <= "100000";
        when "0101110010110" => rgb <= "000000";
        when "0101110010111" => rgb <= "101000";
        when "0101110011000" => rgb <= "101000";
        when "0101110011001" => rgb <= "101000";
        when "0101110011010" => rgb <= "101000";
        when "0101110011011" => rgb <= "101000";
        when "0101110011100" => rgb <= "000000";
        when "0101110011101" => rgb <= "101000";
        when "0101110011110" => rgb <= "101000";
        when "0101110011111" => rgb <= "101000";
        when "0101110100000" => rgb <= "000000";
        when "0101110100100" => rgb <= "000000";
        when "0101110100101" => rgb <= "101000";
        when "0101110100110" => rgb <= "101000";
        when "0101110100111" => rgb <= "101000";
        when "0101110101000" => rgb <= "000000";
        when "0101110101001" => rgb <= "000000";
        when "0101110101010" => rgb <= "001010";
        when "0101110101011" => rgb <= "001010";
        when "0101110101100" => rgb <= "001010";
        when "0101110101101" => rgb <= "000000";
        when "0101110110010" => rgb <= "000000";
        when "0101110110011" => rgb <= "001010";
        when "0101110110100" => rgb <= "001010";
        when "0101110110101" => rgb <= "001010";
        when "0101110110110" => rgb <= "000000";
        when "0101110110111" => rgb <= "100110";
        when "0101110111000" => rgb <= "100110";
        when "0101110111001" => rgb <= "100110";
        when "0101110111010" => rgb <= "100110";
        when "0101110111011" => rgb <= "100110";
        when "0101110111100" => rgb <= "100110";
        when "0101110111101" => rgb <= "100110";
        when "0101110111110" => rgb <= "100110";
        when "0101110111111" => rgb <= "100110";
        when "0101111000000" => rgb <= "100110";
        when "0101111000001" => rgb <= "000000";
        when "0101111000010" => rgb <= "100000";
        when "0101111000011" => rgb <= "100000";
        when "0101111000100" => rgb <= "100000";
        when "0101111000101" => rgb <= "100000";
        when "0101111000110" => rgb <= "100000";
        when "0101111000111" => rgb <= "100000";
        when "0101111001000" => rgb <= "100000";
        when "0101111001001" => rgb <= "000000";
        when "0101111001011" => rgb <= "000000";
        when "0101111001100" => rgb <= "101000";
        when "0101111001101" => rgb <= "000000";
        when "0101111001110" => rgb <= "000000";
        when "0110000000001" => rgb <= "000000";
        when "0110000000010" => rgb <= "100000";
        when "0110000000011" => rgb <= "100000";
        when "0110000000100" => rgb <= "000000";
        when "0110000000101" => rgb <= "000000";
        when "0110000010001" => rgb <= "000000";
        when "0110000010010" => rgb <= "100000";
        when "0110000010011" => rgb <= "100000";
        when "0110000010100" => rgb <= "100000";
        when "0110000010101" => rgb <= "100000";
        when "0110000010110" => rgb <= "000000";
        when "0110000010111" => rgb <= "101000";
        when "0110000011000" => rgb <= "101000";
        when "0110000011001" => rgb <= "101000";
        when "0110000011010" => rgb <= "101000";
        when "0110000011011" => rgb <= "101000";
        when "0110000011100" => rgb <= "000000";
        when "0110000011101" => rgb <= "101000";
        when "0110000011110" => rgb <= "101000";
        when "0110000011111" => rgb <= "101000";
        when "0110000100000" => rgb <= "101000";
        when "0110000100001" => rgb <= "000000";
        when "0110000100100" => rgb <= "000000";
        when "0110000100101" => rgb <= "101000";
        when "0110000100110" => rgb <= "101000";
        when "0110000100111" => rgb <= "101000";
        when "0110000101000" => rgb <= "101000";
        when "0110000101001" => rgb <= "000000";
        when "0110000101010" => rgb <= "001010";
        when "0110000101011" => rgb <= "001010";
        when "0110000101100" => rgb <= "001010";
        when "0110000101101" => rgb <= "001010";
        when "0110000101110" => rgb <= "000000";
        when "0110000110010" => rgb <= "000000";
        when "0110000110011" => rgb <= "001010";
        when "0110000110100" => rgb <= "001010";
        when "0110000110101" => rgb <= "001010";
        when "0110000110110" => rgb <= "000000";
        when "0110000110111" => rgb <= "000000";
        when "0110000111000" => rgb <= "100110";
        when "0110000111001" => rgb <= "100110";
        when "0110000111010" => rgb <= "100110";
        when "0110000111011" => rgb <= "000000";
        when "0110000111100" => rgb <= "000000";
        when "0110000111101" => rgb <= "000000";
        when "0110000111110" => rgb <= "000000";
        when "0110000111111" => rgb <= "000000";
        when "0110001000000" => rgb <= "000000";
        when "0110001000001" => rgb <= "000000";
        when "0110001000010" => rgb <= "100000";
        when "0110001000011" => rgb <= "000000";
        when "0110001000100" => rgb <= "000000";
        when "0110001000101" => rgb <= "000000";
        when "0110001000110" => rgb <= "000000";
        when "0110001000111" => rgb <= "100000";
        when "0110001001000" => rgb <= "100000";
        when "0110001001001" => rgb <= "100000";
        when "0110001001010" => rgb <= "000000";
        when "0110001001011" => rgb <= "000000";
        when "0110001001100" => rgb <= "101000";
        when "0110001001101" => rgb <= "101000";
        when "0110001001110" => rgb <= "000000";
        when "0110010000001" => rgb <= "000000";
        when "0110010000010" => rgb <= "100000";
        when "0110010000011" => rgb <= "100000";
        when "0110010000100" => rgb <= "100000";
        when "0110010000101" => rgb <= "000000";
        when "0110010010000" => rgb <= "000000";
        when "0110010010001" => rgb <= "100000";
        when "0110010010010" => rgb <= "100000";
        when "0110010010011" => rgb <= "100000";
        when "0110010010100" => rgb <= "100000";
        when "0110010010101" => rgb <= "000000";
        when "0110010010110" => rgb <= "101000";
        when "0110010010111" => rgb <= "101000";
        when "0110010011000" => rgb <= "101000";
        when "0110010011001" => rgb <= "000000";
        when "0110010011010" => rgb <= "000000";
        when "0110010011011" => rgb <= "000000";
        when "0110010011100" => rgb <= "101000";
        when "0110010011101" => rgb <= "101000";
        when "0110010011110" => rgb <= "101000";
        when "0110010011111" => rgb <= "101000";
        when "0110010100000" => rgb <= "101000";
        when "0110010100001" => rgb <= "000000";
        when "0110010100101" => rgb <= "000000";
        when "0110010100110" => rgb <= "101000";
        when "0110010100111" => rgb <= "101000";
        when "0110010101000" => rgb <= "101000";
        when "0110010101001" => rgb <= "000000";
        when "0110010101010" => rgb <= "001010";
        when "0110010101011" => rgb <= "001010";
        when "0110010101100" => rgb <= "001010";
        when "0110010101101" => rgb <= "001010";
        when "0110010101110" => rgb <= "001010";
        when "0110010101111" => rgb <= "000000";
        when "0110010110010" => rgb <= "000000";
        when "0110010110011" => rgb <= "001010";
        when "0110010110100" => rgb <= "001010";
        when "0110010110101" => rgb <= "001010";
        when "0110010110110" => rgb <= "001010";
        when "0110010110111" => rgb <= "000000";
        when "0110010111000" => rgb <= "100110";
        when "0110010111001" => rgb <= "100110";
        when "0110010111010" => rgb <= "000000";
        when "0110010111011" => rgb <= "000000";
        when "0110011000000" => rgb <= "000000";
        when "0110011000001" => rgb <= "100000";
        when "0110011000010" => rgb <= "100000";
        when "0110011000011" => rgb <= "000000";
        when "0110011000110" => rgb <= "000000";
        when "0110011000111" => rgb <= "100000";
        when "0110011001000" => rgb <= "100000";
        when "0110011001001" => rgb <= "100000";
        when "0110011001010" => rgb <= "000000";
        when "0110011001011" => rgb <= "000000";
        when "0110011001100" => rgb <= "101000";
        when "0110011001101" => rgb <= "101000";
        when "0110011001110" => rgb <= "000000";
        when "0110100000010" => rgb <= "000000";
        when "0110100000011" => rgb <= "100000";
        when "0110100000100" => rgb <= "100000";
        when "0110100000101" => rgb <= "100000";
        when "0110100000110" => rgb <= "000000";
        when "0110100001111" => rgb <= "000000";
        when "0110100010000" => rgb <= "000000";
        when "0110100010001" => rgb <= "100000";
        when "0110100010010" => rgb <= "100000";
        when "0110100010011" => rgb <= "100000";
        when "0110100010100" => rgb <= "100000";
        when "0110100010101" => rgb <= "000000";
        when "0110100010110" => rgb <= "101000";
        when "0110100010111" => rgb <= "101000";
        when "0110100011000" => rgb <= "101000";
        when "0110100011001" => rgb <= "000000";
        when "0110100011011" => rgb <= "000000";
        when "0110100011100" => rgb <= "101000";
        when "0110100011101" => rgb <= "101000";
        when "0110100011110" => rgb <= "101000";
        when "0110100011111" => rgb <= "101000";
        when "0110100100000" => rgb <= "101000";
        when "0110100100001" => rgb <= "101000";
        when "0110100100010" => rgb <= "000000";
        when "0110100100101" => rgb <= "000000";
        when "0110100100110" => rgb <= "101000";
        when "0110100100111" => rgb <= "101000";
        when "0110100101000" => rgb <= "101000";
        when "0110100101001" => rgb <= "000000";
        when "0110100101010" => rgb <= "001010";
        when "0110100101011" => rgb <= "001010";
        when "0110100101100" => rgb <= "001010";
        when "0110100101101" => rgb <= "001010";
        when "0110100101110" => rgb <= "001010";
        when "0110100101111" => rgb <= "001010";
        when "0110100110000" => rgb <= "000000";
        when "0110100110010" => rgb <= "000000";
        when "0110100110011" => rgb <= "000000";
        when "0110100110100" => rgb <= "001010";
        when "0110100110101" => rgb <= "001010";
        when "0110100110110" => rgb <= "001010";
        when "0110100110111" => rgb <= "000000";
        when "0110100111000" => rgb <= "100110";
        when "0110100111001" => rgb <= "100110";
        when "0110100111010" => rgb <= "000000";
        when "0110101000000" => rgb <= "000000";
        when "0110101000001" => rgb <= "100000";
        when "0110101000010" => rgb <= "100000";
        when "0110101000011" => rgb <= "000000";
        when "0110101000100" => rgb <= "000000";
        when "0110101000101" => rgb <= "000000";
        when "0110101000110" => rgb <= "100000";
        when "0110101000111" => rgb <= "100000";
        when "0110101001000" => rgb <= "100000";
        when "0110101001001" => rgb <= "000000";
        when "0110101001011" => rgb <= "000000";
        when "0110101001100" => rgb <= "000000";
        when "0110101001101" => rgb <= "101000";
        when "0110101001110" => rgb <= "000000";
        when "0110110000010" => rgb <= "000000";
        when "0110110000011" => rgb <= "100000";
        when "0110110000100" => rgb <= "100000";
        when "0110110000101" => rgb <= "100000";
        when "0110110000110" => rgb <= "000000";
        when "0110110001010" => rgb <= "000000";
        when "0110110001011" => rgb <= "000000";
        when "0110110001111" => rgb <= "000000";
        when "0110110010000" => rgb <= "100000";
        when "0110110010001" => rgb <= "100000";
        when "0110110010010" => rgb <= "100000";
        when "0110110010011" => rgb <= "100000";
        when "0110110010100" => rgb <= "000000";
        when "0110110010101" => rgb <= "000000";
        when "0110110010110" => rgb <= "101000";
        when "0110110010111" => rgb <= "101000";
        when "0110110011000" => rgb <= "101000";
        when "0110110011001" => rgb <= "000000";
        when "0110110011011" => rgb <= "000000";
        when "0110110011100" => rgb <= "101000";
        when "0110110011101" => rgb <= "101000";
        when "0110110011110" => rgb <= "101000";
        when "0110110011111" => rgb <= "101000";
        when "0110110100000" => rgb <= "101000";
        when "0110110100001" => rgb <= "101000";
        when "0110110100010" => rgb <= "000000";
        when "0110110100011" => rgb <= "000000";
        when "0110110100101" => rgb <= "000000";
        when "0110110100110" => rgb <= "101000";
        when "0110110100111" => rgb <= "101000";
        when "0110110101000" => rgb <= "101000";
        when "0110110101001" => rgb <= "000000";
        when "0110110101010" => rgb <= "001010";
        when "0110110101011" => rgb <= "001010";
        when "0110110101100" => rgb <= "001010";
        when "0110110101101" => rgb <= "001010";
        when "0110110101110" => rgb <= "001010";
        when "0110110101111" => rgb <= "001010";
        when "0110110110000" => rgb <= "000000";
        when "0110110110001" => rgb <= "000000";
        when "0110110110011" => rgb <= "000000";
        when "0110110110100" => rgb <= "001010";
        when "0110110110101" => rgb <= "001010";
        when "0110110110110" => rgb <= "001010";
        when "0110110110111" => rgb <= "000000";
        when "0110110111000" => rgb <= "100110";
        when "0110110111001" => rgb <= "100110";
        when "0110110111010" => rgb <= "100110";
        when "0110110111011" => rgb <= "000000";
        when "0110110111100" => rgb <= "000000";
        when "0110110111101" => rgb <= "000000";
        when "0110111000000" => rgb <= "000000";
        when "0110111000001" => rgb <= "100000";
        when "0110111000010" => rgb <= "100000";
        when "0110111000011" => rgb <= "100000";
        when "0110111000100" => rgb <= "100000";
        when "0110111000101" => rgb <= "100000";
        when "0110111000110" => rgb <= "100000";
        when "0110111000111" => rgb <= "100000";
        when "0110111001000" => rgb <= "100000";
        when "0110111001001" => rgb <= "000000";
        when "0110111001100" => rgb <= "000000";
        when "0110111001101" => rgb <= "101000";
        when "0110111001110" => rgb <= "000000";
        when "0111000000010" => rgb <= "000000";
        when "0111000000011" => rgb <= "100000";
        when "0111000000100" => rgb <= "100000";
        when "0111000000101" => rgb <= "100000";
        when "0111000000110" => rgb <= "000000";
        when "0111000001000" => rgb <= "000000";
        when "0111000001001" => rgb <= "000000";
        when "0111000001010" => rgb <= "100000";
        when "0111000001011" => rgb <= "000000";
        when "0111000001100" => rgb <= "000000";
        when "0111000001101" => rgb <= "000000";
        when "0111000001110" => rgb <= "000000";
        when "0111000001111" => rgb <= "000000";
        when "0111000010000" => rgb <= "100000";
        when "0111000010001" => rgb <= "100000";
        when "0111000010010" => rgb <= "100000";
        when "0111000010011" => rgb <= "100000";
        when "0111000010100" => rgb <= "000000";
        when "0111000010101" => rgb <= "000000";
        when "0111000010110" => rgb <= "101000";
        when "0111000010111" => rgb <= "101000";
        when "0111000011000" => rgb <= "101000";
        when "0111000011001" => rgb <= "000000";
        when "0111000011011" => rgb <= "000000";
        when "0111000011100" => rgb <= "101000";
        when "0111000011101" => rgb <= "101000";
        when "0111000011110" => rgb <= "101000";
        when "0111000011111" => rgb <= "101000";
        when "0111000100000" => rgb <= "101000";
        when "0111000100001" => rgb <= "101000";
        when "0111000100010" => rgb <= "101000";
        when "0111000100011" => rgb <= "000000";
        when "0111000100101" => rgb <= "000000";
        when "0111000100110" => rgb <= "101000";
        when "0111000100111" => rgb <= "101000";
        when "0111000101000" => rgb <= "101000";
        when "0111000101001" => rgb <= "000000";
        when "0111000101010" => rgb <= "001010";
        when "0111000101011" => rgb <= "001010";
        when "0111000101100" => rgb <= "001010";
        when "0111000101101" => rgb <= "001010";
        when "0111000101110" => rgb <= "001010";
        when "0111000101111" => rgb <= "001010";
        when "0111000110000" => rgb <= "001010";
        when "0111000110001" => rgb <= "000000";
        when "0111000110011" => rgb <= "000000";
        when "0111000110100" => rgb <= "001010";
        when "0111000110101" => rgb <= "001010";
        when "0111000110110" => rgb <= "001010";
        when "0111000110111" => rgb <= "000000";
        when "0111000111000" => rgb <= "100110";
        when "0111000111001" => rgb <= "100110";
        when "0111000111010" => rgb <= "100110";
        when "0111000111011" => rgb <= "100110";
        when "0111000111100" => rgb <= "100110";
        when "0111000111101" => rgb <= "100110";
        when "0111000111110" => rgb <= "000000";
        when "0111001000000" => rgb <= "000000";
        when "0111001000001" => rgb <= "100000";
        when "0111001000010" => rgb <= "100000";
        when "0111001000011" => rgb <= "100000";
        when "0111001000100" => rgb <= "100000";
        when "0111001000101" => rgb <= "100000";
        when "0111001000110" => rgb <= "100000";
        when "0111001000111" => rgb <= "000000";
        when "0111001001000" => rgb <= "000000";
        when "0111001001100" => rgb <= "000000";
        when "0111001001101" => rgb <= "101000";
        when "0111001001110" => rgb <= "000000";
        when "0111010000011" => rgb <= "000000";
        when "0111010000100" => rgb <= "100000";
        when "0111010000101" => rgb <= "100000";
        when "0111010000110" => rgb <= "000000";
        when "0111010000111" => rgb <= "000000";
        when "0111010001000" => rgb <= "000000";
        when "0111010001001" => rgb <= "100000";
        when "0111010001010" => rgb <= "100000";
        when "0111010001011" => rgb <= "100000";
        when "0111010001100" => rgb <= "100000";
        when "0111010001101" => rgb <= "100000";
        when "0111010001110" => rgb <= "100000";
        when "0111010001111" => rgb <= "100000";
        when "0111010010000" => rgb <= "100000";
        when "0111010010001" => rgb <= "100000";
        when "0111010010010" => rgb <= "100000";
        when "0111010010011" => rgb <= "100000";
        when "0111010010100" => rgb <= "000000";
        when "0111010010101" => rgb <= "000000";
        when "0111010010110" => rgb <= "101000";
        when "0111010010111" => rgb <= "101000";
        when "0111010011000" => rgb <= "101000";
        when "0111010011001" => rgb <= "000000";
        when "0111010011011" => rgb <= "000000";
        when "0111010011100" => rgb <= "101000";
        when "0111010011101" => rgb <= "101000";
        when "0111010011110" => rgb <= "101000";
        when "0111010011111" => rgb <= "101000";
        when "0111010100000" => rgb <= "101000";
        when "0111010100001" => rgb <= "101000";
        when "0111010100010" => rgb <= "101000";
        when "0111010100011" => rgb <= "101000";
        when "0111010100100" => rgb <= "000000";
        when "0111010100101" => rgb <= "000000";
        when "0111010100110" => rgb <= "101000";
        when "0111010100111" => rgb <= "101000";
        when "0111010101000" => rgb <= "101000";
        when "0111010101001" => rgb <= "000000";
        when "0111010101010" => rgb <= "001010";
        when "0111010101011" => rgb <= "001010";
        when "0111010101100" => rgb <= "001010";
        when "0111010101101" => rgb <= "000000";
        when "0111010101110" => rgb <= "001010";
        when "0111010101111" => rgb <= "001010";
        when "0111010110000" => rgb <= "001010";
        when "0111010110001" => rgb <= "001010";
        when "0111010110010" => rgb <= "000000";
        when "0111010110011" => rgb <= "000000";
        when "0111010110100" => rgb <= "001010";
        when "0111010110101" => rgb <= "001010";
        when "0111010110110" => rgb <= "001010";
        when "0111010110111" => rgb <= "000000";
        when "0111010111000" => rgb <= "100110";
        when "0111010111001" => rgb <= "100110";
        when "0111010111010" => rgb <= "000000";
        when "0111010111011" => rgb <= "000000";
        when "0111010111100" => rgb <= "000000";
        when "0111010111101" => rgb <= "000000";
        when "0111010111110" => rgb <= "000000";
        when "0111011000000" => rgb <= "000000";
        when "0111011000001" => rgb <= "100000";
        when "0111011000010" => rgb <= "100000";
        when "0111011000011" => rgb <= "100000";
        when "0111011000100" => rgb <= "100000";
        when "0111011000101" => rgb <= "100000";
        when "0111011000110" => rgb <= "100000";
        when "0111011000111" => rgb <= "000000";
        when "0111011001000" => rgb <= "000000";
        when "0111011001100" => rgb <= "000000";
        when "0111011001101" => rgb <= "000000";
        when "0111011001110" => rgb <= "000000";
        when "0111100000011" => rgb <= "000000";
        when "0111100000100" => rgb <= "100000";
        when "0111100000101" => rgb <= "100000";
        when "0111100000110" => rgb <= "100000";
        when "0111100000111" => rgb <= "100000";
        when "0111100001000" => rgb <= "100000";
        when "0111100001001" => rgb <= "100000";
        when "0111100001010" => rgb <= "100000";
        when "0111100001011" => rgb <= "100000";
        when "0111100001100" => rgb <= "100000";
        when "0111100001101" => rgb <= "100000";
        when "0111100001110" => rgb <= "100000";
        when "0111100001111" => rgb <= "100000";
        when "0111100010000" => rgb <= "100000";
        when "0111100010001" => rgb <= "100000";
        when "0111100010010" => rgb <= "100000";
        when "0111100010011" => rgb <= "100000";
        when "0111100010100" => rgb <= "000000";
        when "0111100010101" => rgb <= "000000";
        when "0111100010110" => rgb <= "101000";
        when "0111100010111" => rgb <= "101000";
        when "0111100011000" => rgb <= "101000";
        when "0111100011001" => rgb <= "000000";
        when "0111100011011" => rgb <= "000000";
        when "0111100011100" => rgb <= "101000";
        when "0111100011101" => rgb <= "101000";
        when "0111100011110" => rgb <= "101000";
        when "0111100011111" => rgb <= "101000";
        when "0111100100000" => rgb <= "000000";
        when "0111100100001" => rgb <= "000000";
        when "0111100100010" => rgb <= "101000";
        when "0111100100011" => rgb <= "101000";
        when "0111100100100" => rgb <= "101000";
        when "0111100100101" => rgb <= "000000";
        when "0111100100110" => rgb <= "101000";
        when "0111100100111" => rgb <= "101000";
        when "0111100101000" => rgb <= "101000";
        when "0111100101001" => rgb <= "000000";
        when "0111100101010" => rgb <= "001010";
        when "0111100101011" => rgb <= "001010";
        when "0111100101100" => rgb <= "001010";
        when "0111100101101" => rgb <= "000000";
        when "0111100101110" => rgb <= "000000";
        when "0111100101111" => rgb <= "001010";
        when "0111100110000" => rgb <= "001010";
        when "0111100110001" => rgb <= "001010";
        when "0111100110010" => rgb <= "001010";
        when "0111100110011" => rgb <= "000000";
        when "0111100110100" => rgb <= "001010";
        when "0111100110101" => rgb <= "001010";
        when "0111100110110" => rgb <= "001010";
        when "0111100110111" => rgb <= "000000";
        when "0111100111000" => rgb <= "100110";
        when "0111100111001" => rgb <= "100110";
        when "0111100111010" => rgb <= "000000";
        when "0111101000000" => rgb <= "000000";
        when "0111101000001" => rgb <= "100000";
        when "0111101000010" => rgb <= "100000";
        when "0111101000011" => rgb <= "100000";
        when "0111101000100" => rgb <= "100000";
        when "0111101000101" => rgb <= "100000";
        when "0111101000110" => rgb <= "100000";
        when "0111101000111" => rgb <= "100000";
        when "0111101001000" => rgb <= "100000";
        when "0111101001001" => rgb <= "000000";
        when "0111101001101" => rgb <= "000000";
        when "0111110000011" => rgb <= "000000";
        when "0111110000100" => rgb <= "100000";
        when "0111110000101" => rgb <= "100000";
        when "0111110000110" => rgb <= "100000";
        when "0111110000111" => rgb <= "100000";
        when "0111110001000" => rgb <= "100000";
        when "0111110001001" => rgb <= "100000";
        when "0111110001010" => rgb <= "100000";
        when "0111110001011" => rgb <= "100000";
        when "0111110001100" => rgb <= "100000";
        when "0111110001101" => rgb <= "100000";
        when "0111110001110" => rgb <= "100000";
        when "0111110001111" => rgb <= "100000";
        when "0111110010000" => rgb <= "100000";
        when "0111110010001" => rgb <= "100000";
        when "0111110010010" => rgb <= "100000";
        when "0111110010011" => rgb <= "000000";
        when "0111110010101" => rgb <= "000000";
        when "0111110010110" => rgb <= "101000";
        when "0111110010111" => rgb <= "101000";
        when "0111110011000" => rgb <= "101000";
        when "0111110011001" => rgb <= "000000";
        when "0111110011011" => rgb <= "000000";
        when "0111110011100" => rgb <= "101000";
        when "0111110011101" => rgb <= "101000";
        when "0111110011110" => rgb <= "101000";
        when "0111110011111" => rgb <= "101000";
        when "0111110100000" => rgb <= "000000";
        when "0111110100001" => rgb <= "000000";
        when "0111110100010" => rgb <= "101000";
        when "0111110100011" => rgb <= "101000";
        when "0111110100100" => rgb <= "101000";
        when "0111110100101" => rgb <= "101000";
        when "0111110100110" => rgb <= "101000";
        when "0111110100111" => rgb <= "101000";
        when "0111110101000" => rgb <= "101000";
        when "0111110101001" => rgb <= "000000";
        when "0111110101010" => rgb <= "001010";
        when "0111110101011" => rgb <= "001010";
        when "0111110101100" => rgb <= "001010";
        when "0111110101101" => rgb <= "000000";
        when "0111110101110" => rgb <= "000000";
        when "0111110101111" => rgb <= "001010";
        when "0111110110000" => rgb <= "001010";
        when "0111110110001" => rgb <= "001010";
        when "0111110110010" => rgb <= "001010";
        when "0111110110011" => rgb <= "001010";
        when "0111110110100" => rgb <= "001010";
        when "0111110110101" => rgb <= "001010";
        when "0111110110110" => rgb <= "001010";
        when "0111110110111" => rgb <= "000000";
        when "0111110111000" => rgb <= "100110";
        when "0111110111001" => rgb <= "100110";
        when "0111110111010" => rgb <= "000000";
        when "0111111000000" => rgb <= "000000";
        when "0111111000001" => rgb <= "100000";
        when "0111111000010" => rgb <= "100000";
        when "0111111000011" => rgb <= "100000";
        when "0111111000100" => rgb <= "000000";
        when "0111111000101" => rgb <= "000000";
        when "0111111000110" => rgb <= "100000";
        when "0111111000111" => rgb <= "100000";
        when "0111111001000" => rgb <= "100000";
        when "0111111001001" => rgb <= "000000";
        when "0111111001101" => rgb <= "000000";
        when "1000000000100" => rgb <= "000000";
        when "1000000000101" => rgb <= "100000";
        when "1000000000110" => rgb <= "100000";
        when "1000000000111" => rgb <= "100000";
        when "1000000001000" => rgb <= "100000";
        when "1000000001001" => rgb <= "100000";
        when "1000000001010" => rgb <= "000000";
        when "1000000001011" => rgb <= "000000";
        when "1000000001100" => rgb <= "000000";
        when "1000000001101" => rgb <= "100000";
        when "1000000001110" => rgb <= "100000";
        when "1000000001111" => rgb <= "100000";
        when "1000000010000" => rgb <= "100000";
        when "1000000010001" => rgb <= "100000";
        when "1000000010010" => rgb <= "000000";
        when "1000000010011" => rgb <= "000000";
        when "1000000010101" => rgb <= "000000";
        when "1000000010110" => rgb <= "101000";
        when "1000000010111" => rgb <= "101000";
        when "1000000011000" => rgb <= "101000";
        when "1000000011001" => rgb <= "000000";
        when "1000000011011" => rgb <= "000000";
        when "1000000011100" => rgb <= "101000";
        when "1000000011101" => rgb <= "101000";
        when "1000000011110" => rgb <= "101000";
        when "1000000011111" => rgb <= "101000";
        when "1000000100000" => rgb <= "000000";
        when "1000000100010" => rgb <= "000000";
        when "1000000100011" => rgb <= "000000";
        when "1000000100100" => rgb <= "101000";
        when "1000000100101" => rgb <= "101000";
        when "1000000100110" => rgb <= "101000";
        when "1000000100111" => rgb <= "101000";
        when "1000000101000" => rgb <= "101000";
        when "1000000101001" => rgb <= "000000";
        when "1000000101010" => rgb <= "001010";
        when "1000000101011" => rgb <= "001010";
        when "1000000101100" => rgb <= "001010";
        when "1000000101101" => rgb <= "000000";
        when "1000000101111" => rgb <= "000000";
        when "1000000110000" => rgb <= "000000";
        when "1000000110001" => rgb <= "001010";
        when "1000000110010" => rgb <= "001010";
        when "1000000110011" => rgb <= "001010";
        when "1000000110100" => rgb <= "001010";
        when "1000000110101" => rgb <= "001010";
        when "1000000110110" => rgb <= "001010";
        when "1000000110111" => rgb <= "000000";
        when "1000000111000" => rgb <= "100110";
        when "1000000111001" => rgb <= "100110";
        when "1000000111010" => rgb <= "000000";
        when "1000000111011" => rgb <= "000000";
        when "1000000111100" => rgb <= "000000";
        when "1000000111101" => rgb <= "000000";
        when "1000000111110" => rgb <= "000000";
        when "1000000111111" => rgb <= "000000";
        when "1000001000000" => rgb <= "000000";
        when "1000001000001" => rgb <= "100000";
        when "1000001000010" => rgb <= "100000";
        when "1000001000011" => rgb <= "100000";
        when "1000001000100" => rgb <= "000000";
        when "1000001000110" => rgb <= "000000";
        when "1000001000111" => rgb <= "100000";
        when "1000001001000" => rgb <= "100000";
        when "1000001001001" => rgb <= "100000";
        when "1000001001010" => rgb <= "000000";
        when "1000010000100" => rgb <= "000000";
        when "1000010000101" => rgb <= "100000";
        when "1000010000110" => rgb <= "100000";
        when "1000010000111" => rgb <= "100000";
        when "1000010001000" => rgb <= "100000";
        when "1000010001001" => rgb <= "000000";
        when "1000010001101" => rgb <= "000000";
        when "1000010001110" => rgb <= "100000";
        when "1000010001111" => rgb <= "100000";
        when "1000010010000" => rgb <= "100000";
        when "1000010010001" => rgb <= "100000";
        when "1000010010010" => rgb <= "000000";
        when "1000010010101" => rgb <= "000000";
        when "1000010010110" => rgb <= "101000";
        when "1000010010111" => rgb <= "101000";
        when "1000010011000" => rgb <= "101000";
        when "1000010011001" => rgb <= "000000";
        when "1000010011011" => rgb <= "000000";
        when "1000010011100" => rgb <= "101000";
        when "1000010011101" => rgb <= "101000";
        when "1000010011110" => rgb <= "101000";
        when "1000010011111" => rgb <= "000000";
        when "1000010100000" => rgb <= "000000";
        when "1000010100011" => rgb <= "000000";
        when "1000010100100" => rgb <= "000000";
        when "1000010100101" => rgb <= "101000";
        when "1000010100110" => rgb <= "101000";
        when "1000010100111" => rgb <= "101000";
        when "1000010101000" => rgb <= "101000";
        when "1000010101001" => rgb <= "000000";
        when "1000010101010" => rgb <= "001010";
        when "1000010101011" => rgb <= "001010";
        when "1000010101100" => rgb <= "001010";
        when "1000010101101" => rgb <= "000000";
        when "1000010110000" => rgb <= "000000";
        when "1000010110001" => rgb <= "000000";
        when "1000010110010" => rgb <= "001010";
        when "1000010110011" => rgb <= "001010";
        when "1000010110100" => rgb <= "001010";
        when "1000010110101" => rgb <= "001010";
        when "1000010110110" => rgb <= "001010";
        when "1000010110111" => rgb <= "000000";
        when "1000010111000" => rgb <= "100110";
        when "1000010111001" => rgb <= "100110";
        when "1000010111010" => rgb <= "100110";
        when "1000010111011" => rgb <= "100110";
        when "1000010111100" => rgb <= "100110";
        when "1000010111101" => rgb <= "100110";
        when "1000010111110" => rgb <= "100110";
        when "1000010111111" => rgb <= "100110";
        when "1000011000000" => rgb <= "000000";
        when "1000011000001" => rgb <= "100000";
        when "1000011000010" => rgb <= "100000";
        when "1000011000011" => rgb <= "100000";
        when "1000011000100" => rgb <= "000000";
        when "1000011000110" => rgb <= "000000";
        when "1000011000111" => rgb <= "000000";
        when "1000011001000" => rgb <= "100000";
        when "1000011001001" => rgb <= "100000";
        when "1000011001010" => rgb <= "100000";
        when "1000011001011" => rgb <= "000000";
        when "1000011001100" => rgb <= "000000";
        when "1000011001101" => rgb <= "000000";
        when "1000011001110" => rgb <= "000000";
        when "1000100000101" => rgb <= "000000";
        when "1000100000110" => rgb <= "100000";
        when "1000100000111" => rgb <= "100000";
        when "1000100001000" => rgb <= "100000";
        when "1000100001001" => rgb <= "000000";
        when "1000100001101" => rgb <= "000000";
        when "1000100001110" => rgb <= "100000";
        when "1000100001111" => rgb <= "100000";
        when "1000100010000" => rgb <= "100000";
        when "1000100010001" => rgb <= "000000";
        when "1000100010010" => rgb <= "000000";
        when "1000100010011" => rgb <= "000000";
        when "1000100010100" => rgb <= "000000";
        when "1000100010101" => rgb <= "000000";
        when "1000100010110" => rgb <= "101000";
        when "1000100010111" => rgb <= "101000";
        when "1000100011000" => rgb <= "101000";
        when "1000100011001" => rgb <= "000000";
        when "1000100011010" => rgb <= "000000";
        when "1000100011011" => rgb <= "000000";
        when "1000100011100" => rgb <= "101000";
        when "1000100011101" => rgb <= "101000";
        when "1000100011110" => rgb <= "101000";
        when "1000100011111" => rgb <= "000000";
        when "1000100100100" => rgb <= "000000";
        when "1000100100101" => rgb <= "101000";
        when "1000100100110" => rgb <= "101000";
        when "1000100100111" => rgb <= "101000";
        when "1000100101000" => rgb <= "101000";
        when "1000100101001" => rgb <= "000000";
        when "1000100101010" => rgb <= "001010";
        when "1000100101011" => rgb <= "001010";
        when "1000100101100" => rgb <= "001010";
        when "1000100101101" => rgb <= "000000";
        when "1000100110010" => rgb <= "000000";
        when "1000100110011" => rgb <= "001010";
        when "1000100110100" => rgb <= "001010";
        when "1000100110101" => rgb <= "001010";
        when "1000100110110" => rgb <= "001010";
        when "1000100110111" => rgb <= "000000";
        when "1000100111000" => rgb <= "100110";
        when "1000100111001" => rgb <= "100110";
        when "1000100111010" => rgb <= "100110";
        when "1000100111011" => rgb <= "100110";
        when "1000100111100" => rgb <= "100110";
        when "1000100111101" => rgb <= "100110";
        when "1000100111110" => rgb <= "100110";
        when "1000100111111" => rgb <= "100110";
        when "1000101000000" => rgb <= "100110";
        when "1000101000001" => rgb <= "000000";
        when "1000101000010" => rgb <= "100000";
        when "1000101000011" => rgb <= "100000";
        when "1000101000100" => rgb <= "000000";
        when "1000101000111" => rgb <= "000000";
        when "1000101001000" => rgb <= "100000";
        when "1000101001001" => rgb <= "100000";
        when "1000101001010" => rgb <= "100000";
        when "1000101001011" => rgb <= "000000";
        when "1000101001100" => rgb <= "000000";
        when "1000101001101" => rgb <= "101000";
        when "1000101001110" => rgb <= "000000";
        when "1000110000101" => rgb <= "000000";
        when "1000110000110" => rgb <= "100000";
        when "1000110000111" => rgb <= "100000";
        when "1000110001000" => rgb <= "000000";
        when "1000110001110" => rgb <= "000000";
        when "1000110001111" => rgb <= "000000";
        when "1000110010000" => rgb <= "000000";
        when "1000110010001" => rgb <= "000000";
        when "1000110010010" => rgb <= "101000";
        when "1000110010011" => rgb <= "101000";
        when "1000110010100" => rgb <= "101000";
        when "1000110010101" => rgb <= "101000";
        when "1000110010110" => rgb <= "101000";
        when "1000110010111" => rgb <= "101000";
        when "1000110011000" => rgb <= "101000";
        when "1000110011001" => rgb <= "101000";
        when "1000110011010" => rgb <= "101000";
        when "1000110011011" => rgb <= "101000";
        when "1000110011100" => rgb <= "000000";
        when "1000110011101" => rgb <= "101000";
        when "1000110011110" => rgb <= "101000";
        when "1000110011111" => rgb <= "000000";
        when "1000110100101" => rgb <= "000000";
        when "1000110100110" => rgb <= "101000";
        when "1000110100111" => rgb <= "101000";
        when "1000110101000" => rgb <= "101000";
        when "1000110101001" => rgb <= "000000";
        when "1000110101010" => rgb <= "000000";
        when "1000110101011" => rgb <= "000000";
        when "1000110101100" => rgb <= "001010";
        when "1000110101101" => rgb <= "000000";
        when "1000110110010" => rgb <= "000000";
        when "1000110110011" => rgb <= "000000";
        when "1000110110100" => rgb <= "000000";
        when "1000110110101" => rgb <= "000000";
        when "1000110110110" => rgb <= "000000";
        when "1000110110111" => rgb <= "000000";
        when "1000110111000" => rgb <= "000000";
        when "1000110111001" => rgb <= "000000";
        when "1000110111010" => rgb <= "000000";
        when "1000110111011" => rgb <= "000000";
        when "1000110111100" => rgb <= "000000";
        when "1000110111101" => rgb <= "000000";
        when "1000110111110" => rgb <= "000000";
        when "1000110111111" => rgb <= "000000";
        when "1000111000000" => rgb <= "000000";
        when "1000111000001" => rgb <= "000000";
        when "1000111000010" => rgb <= "000000";
        when "1000111000011" => rgb <= "000000";
        when "1000111000100" => rgb <= "000000";
        when "1000111001000" => rgb <= "000000";
        when "1000111001001" => rgb <= "000000";
        when "1000111001010" => rgb <= "000000";
        when "1000111001011" => rgb <= "000000";
        when "1000111001100" => rgb <= "000000";
        when "1000111001101" => rgb <= "000000";
        when "1000111001110" => rgb <= "000000";
        when "1001000000110" => rgb <= "000000";
        when "1001000000111" => rgb <= "000000";
        when "1001000010000" => rgb <= "000000";
        when "1001000010010" => rgb <= "000000";
        when "1001000010011" => rgb <= "000000";
        when "1001000010100" => rgb <= "000000";
        when "1001000010101" => rgb <= "000000";
        when "1001000010110" => rgb <= "101000";
        when "1001000010111" => rgb <= "101000";
        when "1001000011000" => rgb <= "101000";
        when "1001000011001" => rgb <= "101000";
        when "1001000011010" => rgb <= "000000";
        when "1001000011011" => rgb <= "000000";
        when "1001000011100" => rgb <= "000000";
        when "1001000011101" => rgb <= "000000";
        when "1001000011110" => rgb <= "000000";
        when "1001000011111" => rgb <= "000000";
        when "1001000100110" => rgb <= "000000";
        when "1001000100111" => rgb <= "000000";
        when "1001000101000" => rgb <= "000000";
        when "1001000101001" => rgb <= "000000";
        when "1001000101011" => rgb <= "000000";
        when "1001000101100" => rgb <= "000000";
        when "1001000101101" => rgb <= "000000";
        when "1001010010101" => rgb <= "000000";
        when "1001010010110" => rgb <= "000000";
        when "1001010010111" => rgb <= "000000";
        when "1001010011000" => rgb <= "000000";
        when "1001010011001" => rgb <= "000000";
        when others => rgb <= "001000";
            end case;
   end process;
end Behavioral;