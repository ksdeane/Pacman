library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity start_rom is
   Port (
       x_coord : in std_logic_vector(6 downto 0);
	   y_coord : in std_logic_vector(5 downto 0);
       rgb : out std_logic_vector(5 downto 0)
   );
end start_rom;



architecture Behavioral of start_rom is
signal position : std_logic_vector(12 downto 0);

begin
   process(position)
   begin
	case position is
        when "0100100101111" => rgb <= "000000";
        when "0100100110000" => rgb <= "000000";
        when "0100100110001" => rgb <= "000000";
        when "0100100110010" => rgb <= "000000";
        when "0100110010000" => rgb <= "000000";
        when "0100110010001" => rgb <= "000000";
        when "0100110010010" => rgb <= "000000";
        when "0100110010011" => rgb <= "000000";
        when "0100110010100" => rgb <= "000000";
        when "0100110010101" => rgb <= "000000";
        when "0100110010110" => rgb <= "000000";
        when "0100110010111" => rgb <= "000000";
        when "0100110011000" => rgb <= "000000";
        when "0100110011001" => rgb <= "000000";
        when "0100110011010" => rgb <= "000000";
        when "0100110011011" => rgb <= "000000";
        when "0100110011100" => rgb <= "000000";
        when "0100110011101" => rgb <= "000000";
        when "0100110011110" => rgb <= "000000";
        when "0100110100001" => rgb <= "000000";
        when "0100110100010" => rgb <= "000000";
        when "0100110100011" => rgb <= "000000";
        when "0100110100100" => rgb <= "000000";
        when "0100110100101" => rgb <= "000000";
        when "0100110100110" => rgb <= "000000";
        when "0100110100111" => rgb <= "000000";
        when "0100110101000" => rgb <= "000000";
        when "0100110101001" => rgb <= "000000";
        when "0100110101100" => rgb <= "000000";
        when "0100110101101" => rgb <= "000000";
        when "0100110101110" => rgb <= "000000";
        when "0100110101111" => rgb <= "100110";
        when "0100110110000" => rgb <= "100110";
        when "0100110110001" => rgb <= "100110";
        when "0100110110010" => rgb <= "100110";
        when "0100110110011" => rgb <= "000000";
        when "0100110110100" => rgb <= "000000";
        when "0100110110101" => rgb <= "000000";
        when "0100110110110" => rgb <= "000000";
        when "0100110110111" => rgb <= "000000";
        when "0100110111000" => rgb <= "000000";
        when "0100110111001" => rgb <= "000000";
        when "0100110111010" => rgb <= "000000";
        when "0100110111011" => rgb <= "000000";
        when "0100110111100" => rgb <= "000000";
        when "0100110111101" => rgb <= "000000";
        when "0100110111110" => rgb <= "000000";
        when "0100110111111" => rgb <= "000000";
        when "0100111000000" => rgb <= "000000";
        when "0100111000001" => rgb <= "000000";
        when "0100111000010" => rgb <= "000000";
        when "0100111000011" => rgb <= "000000";
        when "0100111000100" => rgb <= "000000";
        when "0100111000101" => rgb <= "000000";
        when "0101000001100" => rgb <= "000000";
        when "0101000001101" => rgb <= "000000";
        when "0101000001110" => rgb <= "000000";
        when "0101000001111" => rgb <= "000000";
        when "0101000010000" => rgb <= "000000";
        when "0101000010001" => rgb <= "000000";
        when "0101000010010" => rgb <= "101000";
        when "0101000010011" => rgb <= "101000";
        when "0101000010100" => rgb <= "101000";
        when "0101000010101" => rgb <= "101000";
        when "0101000010110" => rgb <= "101000";
        when "0101000010111" => rgb <= "101000";
        when "0101000011000" => rgb <= "101000";
        when "0101000011001" => rgb <= "101000";
        when "0101000011010" => rgb <= "101000";
        when "0101000011011" => rgb <= "101000";
        when "0101000011100" => rgb <= "101000";
        when "0101000011101" => rgb <= "101000";
        when "0101000011110" => rgb <= "101000";
        when "0101000011111" => rgb <= "000000";
        when "0101000100000" => rgb <= "000000";
        when "0101000100001" => rgb <= "000000";
        when "0101000100010" => rgb <= "001010";
        when "0101000100011" => rgb <= "001010";
        when "0101000100100" => rgb <= "001010";
        when "0101000100101" => rgb <= "001010";
        when "0101000100110" => rgb <= "001010";
        when "0101000100111" => rgb <= "001010";
        when "0101000101000" => rgb <= "001010";
        when "0101000101001" => rgb <= "001010";
        when "0101000101010" => rgb <= "000000";
        when "0101000101100" => rgb <= "000000";
        when "0101000101101" => rgb <= "100110";
        when "0101000101110" => rgb <= "100110";
        when "0101000101111" => rgb <= "100110";
        when "0101000110000" => rgb <= "100110";
        when "0101000110001" => rgb <= "100110";
        when "0101000110010" => rgb <= "100110";
        when "0101000110011" => rgb <= "100110";
        when "0101000110100" => rgb <= "100110";
        when "0101000110101" => rgb <= "100110";
        when "0101000110110" => rgb <= "000000";
        when "0101000110111" => rgb <= "000000";
        when "0101000111000" => rgb <= "101000";
        when "0101000111001" => rgb <= "101000";
        when "0101000111010" => rgb <= "101000";
        when "0101000111011" => rgb <= "101000";
        when "0101000111100" => rgb <= "101000";
        when "0101000111101" => rgb <= "101000";
        when "0101000111110" => rgb <= "101000";
        when "0101000111111" => rgb <= "101000";
        when "0101001000000" => rgb <= "101000";
        when "0101001000001" => rgb <= "101000";
        when "0101001000010" => rgb <= "101000";
        when "0101001000011" => rgb <= "101000";
        when "0101001000100" => rgb <= "101000";
        when "0101001000101" => rgb <= "000000";
        when "0101010001011" => rgb <= "000000";
        when "0101010001100" => rgb <= "000000";
        when "0101010001101" => rgb <= "100000";
        when "0101010001110" => rgb <= "100000";
        when "0101010001111" => rgb <= "100000";
        when "0101010010000" => rgb <= "100000";
        when "0101010010001" => rgb <= "000000";
        when "0101010010010" => rgb <= "000000";
        when "0101010010011" => rgb <= "101000";
        when "0101010010100" => rgb <= "101000";
        when "0101010010101" => rgb <= "101000";
        when "0101010010110" => rgb <= "101000";
        when "0101010010111" => rgb <= "101000";
        when "0101010011000" => rgb <= "101000";
        when "0101010011001" => rgb <= "101000";
        when "0101010011010" => rgb <= "101000";
        when "0101010011011" => rgb <= "101000";
        when "0101010011100" => rgb <= "101000";
        when "0101010011101" => rgb <= "101000";
        when "0101010011110" => rgb <= "101000";
        when "0101010011111" => rgb <= "101000";
        when "0101010100000" => rgb <= "000000";
        when "0101010100001" => rgb <= "001010";
        when "0101010100010" => rgb <= "001010";
        when "0101010100011" => rgb <= "001010";
        when "0101010100100" => rgb <= "001010";
        when "0101010100101" => rgb <= "001010";
        when "0101010100110" => rgb <= "001010";
        when "0101010100111" => rgb <= "001010";
        when "0101010101000" => rgb <= "001010";
        when "0101010101001" => rgb <= "001010";
        when "0101010101010" => rgb <= "001010";
        when "0101010101011" => rgb <= "000000";
        when "0101010101100" => rgb <= "000000";
        when "0101010101101" => rgb <= "100110";
        when "0101010101110" => rgb <= "100110";
        when "0101010101111" => rgb <= "100110";
        when "0101010110000" => rgb <= "100110";
        when "0101010110001" => rgb <= "100110";
        when "0101010110010" => rgb <= "100110";
        when "0101010110011" => rgb <= "100110";
        when "0101010110100" => rgb <= "100110";
        when "0101010110101" => rgb <= "100110";
        when "0101010110110" => rgb <= "100110";
        when "0101010110111" => rgb <= "000000";
        when "0101010111000" => rgb <= "000000";
        when "0101010111001" => rgb <= "101000";
        when "0101010111010" => rgb <= "101000";
        when "0101010111011" => rgb <= "101000";
        when "0101010111100" => rgb <= "101000";
        when "0101010111101" => rgb <= "101000";
        when "0101010111110" => rgb <= "101000";
        when "0101010111111" => rgb <= "101000";
        when "0101011000000" => rgb <= "101000";
        when "0101011000001" => rgb <= "101000";
        when "0101011000010" => rgb <= "101000";
        when "0101011000011" => rgb <= "101000";
        when "0101011000100" => rgb <= "101000";
        when "0101011000101" => rgb <= "000000";
        when "0101100001010" => rgb <= "000000";
        when "0101100001011" => rgb <= "100000";
        when "0101100001100" => rgb <= "100000";
        when "0101100001101" => rgb <= "100000";
        when "0101100001110" => rgb <= "100000";
        when "0101100001111" => rgb <= "100000";
        when "0101100010000" => rgb <= "100000";
        when "0101100010001" => rgb <= "100000";
        when "0101100010010" => rgb <= "000000";
        when "0101100010011" => rgb <= "101000";
        when "0101100010100" => rgb <= "101000";
        when "0101100010101" => rgb <= "101000";
        when "0101100010110" => rgb <= "101000";
        when "0101100010111" => rgb <= "101000";
        when "0101100011000" => rgb <= "101000";
        when "0101100011001" => rgb <= "101000";
        when "0101100011010" => rgb <= "101000";
        when "0101100011011" => rgb <= "101000";
        when "0101100011100" => rgb <= "101000";
        when "0101100011101" => rgb <= "101000";
        when "0101100011110" => rgb <= "101000";
        when "0101100011111" => rgb <= "000000";
        when "0101100100000" => rgb <= "000000";
        when "0101100100001" => rgb <= "001010";
        when "0101100100010" => rgb <= "001010";
        when "0101100100011" => rgb <= "001010";
        when "0101100100100" => rgb <= "001010";
        when "0101100100101" => rgb <= "001010";
        when "0101100100110" => rgb <= "001010";
        when "0101100100111" => rgb <= "001010";
        when "0101100101000" => rgb <= "001010";
        when "0101100101001" => rgb <= "001010";
        when "0101100101010" => rgb <= "001010";
        when "0101100101011" => rgb <= "000000";
        when "0101100101100" => rgb <= "000000";
        when "0101100101101" => rgb <= "100110";
        when "0101100101110" => rgb <= "100110";
        when "0101100101111" => rgb <= "100110";
        when "0101100110000" => rgb <= "100110";
        when "0101100110001" => rgb <= "100110";
        when "0101100110010" => rgb <= "100110";
        when "0101100110011" => rgb <= "100110";
        when "0101100110100" => rgb <= "100110";
        when "0101100110101" => rgb <= "100110";
        when "0101100110110" => rgb <= "100110";
        when "0101100110111" => rgb <= "100110";
        when "0101100111000" => rgb <= "000000";
        when "0101100111001" => rgb <= "000000";
        when "0101100111010" => rgb <= "000000";
        when "0101100111011" => rgb <= "000000";
        when "0101100111100" => rgb <= "101000";
        when "0101100111101" => rgb <= "101000";
        when "0101100111110" => rgb <= "101000";
        when "0101100111111" => rgb <= "101000";
        when "0101101000000" => rgb <= "000000";
        when "0101101000001" => rgb <= "000000";
        when "0101101000010" => rgb <= "000000";
        when "0101101000011" => rgb <= "000000";
        when "0101101000100" => rgb <= "000000";
        when "0101101000101" => rgb <= "000000";
        when "0101110001001" => rgb <= "000000";
        when "0101110001010" => rgb <= "100000";
        when "0101110001011" => rgb <= "100000";
        when "0101110001100" => rgb <= "100000";
        when "0101110001101" => rgb <= "100000";
        when "0101110001110" => rgb <= "100000";
        when "0101110001111" => rgb <= "100000";
        when "0101110010000" => rgb <= "000000";
        when "0101110010001" => rgb <= "000000";
        when "0101110010010" => rgb <= "000000";
        when "0101110010011" => rgb <= "000000";
        when "0101110010100" => rgb <= "000000";
        when "0101110010101" => rgb <= "000000";
        when "0101110010110" => rgb <= "000000";
        when "0101110010111" => rgb <= "000000";
        when "0101110011000" => rgb <= "101000";
        when "0101110011001" => rgb <= "101000";
        when "0101110011010" => rgb <= "101000";
        when "0101110011011" => rgb <= "000000";
        when "0101110011100" => rgb <= "000000";
        when "0101110011101" => rgb <= "000000";
        when "0101110011110" => rgb <= "000000";
        when "0101110011111" => rgb <= "000000";
        when "0101110100000" => rgb <= "001010";
        when "0101110100001" => rgb <= "001010";
        when "0101110100010" => rgb <= "000000";
        when "0101110100011" => rgb <= "000000";
        when "0101110100100" => rgb <= "000000";
        when "0101110100101" => rgb <= "000000";
        when "0101110100110" => rgb <= "001010";
        when "0101110100111" => rgb <= "000000";
        when "0101110101000" => rgb <= "000000";
        when "0101110101001" => rgb <= "000000";
        when "0101110101010" => rgb <= "000000";
        when "0101110101011" => rgb <= "001010";
        when "0101110101100" => rgb <= "000000";
        when "0101110101101" => rgb <= "000000";
        when "0101110101110" => rgb <= "100110";
        when "0101110101111" => rgb <= "100110";
        when "0101110110000" => rgb <= "000000";
        when "0101110110001" => rgb <= "000000";
        when "0101110110010" => rgb <= "000000";
        when "0101110110011" => rgb <= "000000";
        when "0101110110100" => rgb <= "100110";
        when "0101110110101" => rgb <= "100110";
        when "0101110110110" => rgb <= "100110";
        when "0101110110111" => rgb <= "100110";
        when "0101110111000" => rgb <= "100110";
        when "0101110111001" => rgb <= "000000";
        when "0101110111100" => rgb <= "000000";
        when "0101110111101" => rgb <= "101000";
        when "0101110111110" => rgb <= "101000";
        when "0101110111111" => rgb <= "101000";
        when "0101111000000" => rgb <= "000000";
        when "0110000001001" => rgb <= "000000";
        when "0110000001010" => rgb <= "100000";
        when "0110000001011" => rgb <= "100000";
        when "0110000001100" => rgb <= "100000";
        when "0110000001101" => rgb <= "100000";
        when "0110000001110" => rgb <= "100000";
        when "0110000001111" => rgb <= "000000";
        when "0110000010111" => rgb <= "000000";
        when "0110000011000" => rgb <= "101000";
        when "0110000011001" => rgb <= "101000";
        when "0110000011010" => rgb <= "101000";
        when "0110000011011" => rgb <= "000000";
        when "0110000011110" => rgb <= "000000";
        when "0110000011111" => rgb <= "000000";
        when "0110000100000" => rgb <= "001010";
        when "0110000100001" => rgb <= "001010";
        when "0110000100010" => rgb <= "000000";
        when "0110000100011" => rgb <= "000000";
        when "0110000100100" => rgb <= "101010";
        when "0110000100101" => rgb <= "000000";
        when "0110000100110" => rgb <= "001010";
        when "0110000100111" => rgb <= "000000";
        when "0110000101000" => rgb <= "000000";
        when "0110000101001" => rgb <= "101010";
        when "0110000101010" => rgb <= "000000";
        when "0110000101011" => rgb <= "001010";
        when "0110000101100" => rgb <= "001010";
        when "0110000101101" => rgb <= "000000";
        when "0110000101110" => rgb <= "100110";
        when "0110000101111" => rgb <= "100110";
        when "0110000110000" => rgb <= "000000";
        when "0110000110011" => rgb <= "000000";
        when "0110000110100" => rgb <= "100110";
        when "0110000110101" => rgb <= "100110";
        when "0110000110110" => rgb <= "100110";
        when "0110000110111" => rgb <= "100110";
        when "0110000111000" => rgb <= "100110";
        when "0110000111001" => rgb <= "000000";
        when "0110000111100" => rgb <= "000000";
        when "0110000111101" => rgb <= "101000";
        when "0110000111110" => rgb <= "101000";
        when "0110000111111" => rgb <= "101000";
        when "0110001000000" => rgb <= "000000";
        when "0110010001001" => rgb <= "000000";
        when "0110010001010" => rgb <= "100000";
        when "0110010001011" => rgb <= "100000";
        when "0110010001100" => rgb <= "100000";
        when "0110010001101" => rgb <= "100000";
        when "0110010001110" => rgb <= "100000";
        when "0110010001111" => rgb <= "000000";
        when "0110010010111" => rgb <= "000000";
        when "0110010011000" => rgb <= "101000";
        when "0110010011001" => rgb <= "101000";
        when "0110010011010" => rgb <= "101000";
        when "0110010011011" => rgb <= "000000";
        when "0110010011110" => rgb <= "000000";
        when "0110010011111" => rgb <= "001010";
        when "0110010100000" => rgb <= "001010";
        when "0110010100001" => rgb <= "001010";
        when "0110010100010" => rgb <= "000000";
        when "0110010100011" => rgb <= "000000";
        when "0110010100100" => rgb <= "101010";
        when "0110010100101" => rgb <= "000000";
        when "0110010100110" => rgb <= "001010";
        when "0110010100111" => rgb <= "000000";
        when "0110010101000" => rgb <= "000000";
        when "0110010101001" => rgb <= "101010";
        when "0110010101010" => rgb <= "000000";
        when "0110010101011" => rgb <= "001010";
        when "0110010101100" => rgb <= "001010";
        when "0110010101101" => rgb <= "000000";
        when "0110010101110" => rgb <= "100110";
        when "0110010101111" => rgb <= "100110";
        when "0110010110000" => rgb <= "000000";
        when "0110010110001" => rgb <= "000000";
        when "0110010110010" => rgb <= "000000";
        when "0110010110011" => rgb <= "000000";
        when "0110010110100" => rgb <= "100110";
        when "0110010110101" => rgb <= "100110";
        when "0110010110110" => rgb <= "100110";
        when "0110010110111" => rgb <= "100110";
        when "0110010111000" => rgb <= "100110";
        when "0110010111001" => rgb <= "000000";
        when "0110010111100" => rgb <= "000000";
        when "0110010111101" => rgb <= "101000";
        when "0110010111110" => rgb <= "101000";
        when "0110010111111" => rgb <= "101000";
        when "0110011000000" => rgb <= "000000";
        when "0110100001001" => rgb <= "000000";
        when "0110100001010" => rgb <= "100000";
        when "0110100001011" => rgb <= "100000";
        when "0110100001100" => rgb <= "100000";
        when "0110100001101" => rgb <= "100000";
        when "0110100001110" => rgb <= "100000";
        when "0110100001111" => rgb <= "100000";
        when "0110100010000" => rgb <= "000000";
        when "0110100010111" => rgb <= "000000";
        when "0110100011000" => rgb <= "101000";
        when "0110100011001" => rgb <= "101000";
        when "0110100011010" => rgb <= "101000";
        when "0110100011011" => rgb <= "000000";
        when "0110100011110" => rgb <= "000000";
        when "0110100011111" => rgb <= "001010";
        when "0110100100000" => rgb <= "001010";
        when "0110100100001" => rgb <= "001010";
        when "0110100100010" => rgb <= "000000";
        when "0110100100011" => rgb <= "101010";
        when "0110100100100" => rgb <= "101010";
        when "0110100100101" => rgb <= "000000";
        when "0110100100110" => rgb <= "001010";
        when "0110100100111" => rgb <= "000000";
        when "0110100101000" => rgb <= "101010";
        when "0110100101001" => rgb <= "101010";
        when "0110100101010" => rgb <= "000000";
        when "0110100101011" => rgb <= "001010";
        when "0110100101100" => rgb <= "001010";
        when "0110100101101" => rgb <= "000000";
        when "0110100101110" => rgb <= "100110";
        when "0110100101111" => rgb <= "100110";
        when "0110100110000" => rgb <= "100110";
        when "0110100110001" => rgb <= "100110";
        when "0110100110010" => rgb <= "100110";
        when "0110100110011" => rgb <= "100110";
        when "0110100110100" => rgb <= "100110";
        when "0110100110101" => rgb <= "100110";
        when "0110100110110" => rgb <= "100110";
        when "0110100110111" => rgb <= "100110";
        when "0110100111000" => rgb <= "100110";
        when "0110100111001" => rgb <= "000000";
        when "0110100111100" => rgb <= "000000";
        when "0110100111101" => rgb <= "101000";
        when "0110100111110" => rgb <= "101000";
        when "0110100111111" => rgb <= "101000";
        when "0110101000000" => rgb <= "000000";
        when "0110110001010" => rgb <= "000000";
        when "0110110001011" => rgb <= "000000";
        when "0110110001100" => rgb <= "100000";
        when "0110110001101" => rgb <= "100000";
        when "0110110001110" => rgb <= "100000";
        when "0110110001111" => rgb <= "100000";
        when "0110110010000" => rgb <= "100000";
        when "0110110010001" => rgb <= "000000";
        when "0110110010010" => rgb <= "000000";
        when "0110110010111" => rgb <= "000000";
        when "0110110011000" => rgb <= "101000";
        when "0110110011001" => rgb <= "101000";
        when "0110110011010" => rgb <= "101000";
        when "0110110011011" => rgb <= "000000";
        when "0110110011110" => rgb <= "000000";
        when "0110110011111" => rgb <= "001010";
        when "0110110100000" => rgb <= "001010";
        when "0110110100001" => rgb <= "001010";
        when "0110110100010" => rgb <= "000000";
        when "0110110100011" => rgb <= "000000";
        when "0110110100100" => rgb <= "000000";
        when "0110110100101" => rgb <= "000000";
        when "0110110100110" => rgb <= "001010";
        when "0110110100111" => rgb <= "000000";
        when "0110110101000" => rgb <= "000000";
        when "0110110101001" => rgb <= "000000";
        when "0110110101010" => rgb <= "000000";
        when "0110110101011" => rgb <= "001010";
        when "0110110101100" => rgb <= "001010";
        when "0110110101101" => rgb <= "000000";
        when "0110110101110" => rgb <= "100110";
        when "0110110101111" => rgb <= "100110";
        when "0110110110000" => rgb <= "100110";
        when "0110110110001" => rgb <= "100110";
        when "0110110110010" => rgb <= "100110";
        when "0110110110011" => rgb <= "100110";
        when "0110110110100" => rgb <= "100110";
        when "0110110110101" => rgb <= "100110";
        when "0110110110110" => rgb <= "100110";
        when "0110110110111" => rgb <= "100110";
        when "0110110111000" => rgb <= "000000";
        when "0110110111100" => rgb <= "000000";
        when "0110110111101" => rgb <= "101000";
        when "0110110111110" => rgb <= "101000";
        when "0110110111111" => rgb <= "101000";
        when "0110111000000" => rgb <= "000000";
        when "0111000001011" => rgb <= "000000";
        when "0111000001100" => rgb <= "000000";
        when "0111000001101" => rgb <= "000000";
        when "0111000001110" => rgb <= "100000";
        when "0111000001111" => rgb <= "100000";
        when "0111000010000" => rgb <= "100000";
        when "0111000010001" => rgb <= "100000";
        when "0111000010010" => rgb <= "000000";
        when "0111000010111" => rgb <= "000000";
        when "0111000011000" => rgb <= "101000";
        when "0111000011001" => rgb <= "101000";
        when "0111000011010" => rgb <= "101000";
        when "0111000011011" => rgb <= "000000";
        when "0111000011110" => rgb <= "000000";
        when "0111000011111" => rgb <= "001010";
        when "0111000100000" => rgb <= "001010";
        when "0111000100001" => rgb <= "001010";
        when "0111000100010" => rgb <= "001010";
        when "0111000100011" => rgb <= "001010";
        when "0111000100100" => rgb <= "001010";
        when "0111000100101" => rgb <= "001010";
        when "0111000100110" => rgb <= "001010";
        when "0111000100111" => rgb <= "001010";
        when "0111000101000" => rgb <= "001010";
        when "0111000101001" => rgb <= "001010";
        when "0111000101010" => rgb <= "001010";
        when "0111000101011" => rgb <= "001010";
        when "0111000101100" => rgb <= "001010";
        when "0111000101101" => rgb <= "000000";
        when "0111000101110" => rgb <= "100110";
        when "0111000101111" => rgb <= "100110";
        when "0111000110000" => rgb <= "100110";
        when "0111000110001" => rgb <= "100110";
        when "0111000110010" => rgb <= "100110";
        when "0111000110011" => rgb <= "100110";
        when "0111000110100" => rgb <= "100110";
        when "0111000110101" => rgb <= "100110";
        when "0111000110110" => rgb <= "100110";
        when "0111000110111" => rgb <= "000000";
        when "0111000111000" => rgb <= "000000";
        when "0111000111100" => rgb <= "000000";
        when "0111000111101" => rgb <= "101000";
        when "0111000111110" => rgb <= "101000";
        when "0111000111111" => rgb <= "101000";
        when "0111001000000" => rgb <= "000000";
        when "0111010001110" => rgb <= "000000";
        when "0111010001111" => rgb <= "100000";
        when "0111010010000" => rgb <= "100000";
        when "0111010010001" => rgb <= "100000";
        when "0111010010010" => rgb <= "100000";
        when "0111010010011" => rgb <= "000000";
        when "0111010010111" => rgb <= "000000";
        when "0111010011000" => rgb <= "101000";
        when "0111010011001" => rgb <= "101000";
        when "0111010011010" => rgb <= "101000";
        when "0111010011011" => rgb <= "000000";
        when "0111010011110" => rgb <= "000000";
        when "0111010011111" => rgb <= "001010";
        when "0111010100000" => rgb <= "001010";
        when "0111010100001" => rgb <= "001010";
        when "0111010100010" => rgb <= "001010";
        when "0111010100011" => rgb <= "001010";
        when "0111010100100" => rgb <= "001010";
        when "0111010100101" => rgb <= "001010";
        when "0111010100110" => rgb <= "001010";
        when "0111010100111" => rgb <= "001010";
        when "0111010101000" => rgb <= "001010";
        when "0111010101001" => rgb <= "001010";
        when "0111010101010" => rgb <= "001010";
        when "0111010101011" => rgb <= "001010";
        when "0111010101100" => rgb <= "001010";
        when "0111010101101" => rgb <= "000000";
        when "0111010101110" => rgb <= "100110";
        when "0111010101111" => rgb <= "100110";
        when "0111010110000" => rgb <= "100110";
        when "0111010110001" => rgb <= "100110";
        when "0111010110010" => rgb <= "100110";
        when "0111010110011" => rgb <= "100110";
        when "0111010110100" => rgb <= "100110";
        when "0111010110101" => rgb <= "000000";
        when "0111010110110" => rgb <= "000000";
        when "0111010111100" => rgb <= "000000";
        when "0111010111101" => rgb <= "101000";
        when "0111010111110" => rgb <= "101000";
        when "0111010111111" => rgb <= "101000";
        when "0111011000000" => rgb <= "000000";
        when "0111100001111" => rgb <= "000000";
        when "0111100010000" => rgb <= "100000";
        when "0111100010001" => rgb <= "100000";
        when "0111100010010" => rgb <= "100000";
        when "0111100010011" => rgb <= "100000";
        when "0111100010100" => rgb <= "000000";
        when "0111100010111" => rgb <= "000000";
        when "0111100011000" => rgb <= "101000";
        when "0111100011001" => rgb <= "101000";
        when "0111100011010" => rgb <= "101000";
        when "0111100011011" => rgb <= "000000";
        when "0111100011110" => rgb <= "000000";
        when "0111100011111" => rgb <= "001010";
        when "0111100100000" => rgb <= "001010";
        when "0111100100001" => rgb <= "001010";
        when "0111100100010" => rgb <= "001010";
        when "0111100100011" => rgb <= "001010";
        when "0111100100100" => rgb <= "001010";
        when "0111100100101" => rgb <= "001010";
        when "0111100100110" => rgb <= "001010";
        when "0111100100111" => rgb <= "001010";
        when "0111100101000" => rgb <= "001010";
        when "0111100101001" => rgb <= "001010";
        when "0111100101010" => rgb <= "001010";
        when "0111100101011" => rgb <= "001010";
        when "0111100101100" => rgb <= "001010";
        when "0111100101101" => rgb <= "000000";
        when "0111100101110" => rgb <= "100110";
        when "0111100101111" => rgb <= "100110";
        when "0111100110000" => rgb <= "100110";
        when "0111100110001" => rgb <= "000000";
        when "0111100110010" => rgb <= "000000";
        when "0111100110011" => rgb <= "100110";
        when "0111100110100" => rgb <= "100110";
        when "0111100110101" => rgb <= "100110";
        when "0111100110110" => rgb <= "000000";
        when "0111100110111" => rgb <= "000000";
        when "0111100111100" => rgb <= "000000";
        when "0111100111101" => rgb <= "101000";
        when "0111100111110" => rgb <= "101000";
        when "0111100111111" => rgb <= "101000";
        when "0111101000000" => rgb <= "000000";
        when "0111110001111" => rgb <= "000000";
        when "0111110010000" => rgb <= "100000";
        when "0111110010001" => rgb <= "100000";
        when "0111110010010" => rgb <= "100000";
        when "0111110010011" => rgb <= "100000";
        when "0111110010100" => rgb <= "000000";
        when "0111110010111" => rgb <= "000000";
        when "0111110011000" => rgb <= "101000";
        when "0111110011001" => rgb <= "101000";
        when "0111110011010" => rgb <= "101000";
        when "0111110011011" => rgb <= "000000";
        when "0111110011110" => rgb <= "000000";
        when "0111110011111" => rgb <= "001010";
        when "0111110100000" => rgb <= "001010";
        when "0111110100001" => rgb <= "001010";
        when "0111110100010" => rgb <= "001010";
        when "0111110100011" => rgb <= "001010";
        when "0111110100100" => rgb <= "001010";
        when "0111110100101" => rgb <= "001010";
        when "0111110100110" => rgb <= "001010";
        when "0111110100111" => rgb <= "001010";
        when "0111110101000" => rgb <= "001010";
        when "0111110101001" => rgb <= "001010";
        when "0111110101010" => rgb <= "001010";
        when "0111110101011" => rgb <= "001010";
        when "0111110101100" => rgb <= "001010";
        when "0111110101101" => rgb <= "000000";
        when "0111110101110" => rgb <= "100110";
        when "0111110101111" => rgb <= "100110";
        when "0111110110000" => rgb <= "100110";
        when "0111110110001" => rgb <= "000000";
        when "0111110110010" => rgb <= "000000";
        when "0111110110011" => rgb <= "000000";
        when "0111110110100" => rgb <= "100110";
        when "0111110110101" => rgb <= "100110";
        when "0111110110110" => rgb <= "000000";
        when "0111110110111" => rgb <= "000000";
        when "0111110111100" => rgb <= "000000";
        when "0111110111101" => rgb <= "101000";
        when "0111110111110" => rgb <= "101000";
        when "0111110111111" => rgb <= "101000";
        when "0111111000000" => rgb <= "000000";
        when "1000000000111" => rgb <= "000000";
        when "1000000001000" => rgb <= "000000";
        when "1000000001001" => rgb <= "000000";
        when "1000000001111" => rgb <= "000000";
        when "1000000010000" => rgb <= "000000";
        when "1000000010001" => rgb <= "100000";
        when "1000000010010" => rgb <= "100000";
        when "1000000010011" => rgb <= "100000";
        when "1000000010100" => rgb <= "000000";
        when "1000000010111" => rgb <= "000000";
        when "1000000011000" => rgb <= "101000";
        when "1000000011001" => rgb <= "101000";
        when "1000000011010" => rgb <= "101000";
        when "1000000011011" => rgb <= "000000";
        when "1000000011110" => rgb <= "000000";
        when "1000000011111" => rgb <= "001010";
        when "1000000100000" => rgb <= "001010";
        when "1000000100001" => rgb <= "001010";
        when "1000000100010" => rgb <= "001010";
        when "1000000100011" => rgb <= "001010";
        when "1000000100100" => rgb <= "001010";
        when "1000000100101" => rgb <= "001010";
        when "1000000100110" => rgb <= "001010";
        when "1000000100111" => rgb <= "001010";
        when "1000000101000" => rgb <= "001010";
        when "1000000101001" => rgb <= "001010";
        when "1000000101010" => rgb <= "001010";
        when "1000000101011" => rgb <= "001010";
        when "1000000101100" => rgb <= "001010";
        when "1000000101101" => rgb <= "000000";
        when "1000000101110" => rgb <= "100110";
        when "1000000101111" => rgb <= "100110";
        when "1000000110000" => rgb <= "100110";
        when "1000000110001" => rgb <= "000000";
        when "1000000110011" => rgb <= "000000";
        when "1000000110100" => rgb <= "000000";
        when "1000000110101" => rgb <= "100110";
        when "1000000110110" => rgb <= "100110";
        when "1000000110111" => rgb <= "100110";
        when "1000000111000" => rgb <= "000000";
        when "1000000111100" => rgb <= "000000";
        when "1000000111101" => rgb <= "101000";
        when "1000000111110" => rgb <= "101000";
        when "1000000111111" => rgb <= "101000";
        when "1000001000000" => rgb <= "000000";
        when "1000010000110" => rgb <= "000000";
        when "1000010000111" => rgb <= "100000";
        when "1000010001000" => rgb <= "100000";
        when "1000010001001" => rgb <= "100000";
        when "1000010001010" => rgb <= "000000";
        when "1000010001011" => rgb <= "000000";
        when "1000010001110" => rgb <= "000000";
        when "1000010001111" => rgb <= "000000";
        when "1000010010000" => rgb <= "100000";
        when "1000010010001" => rgb <= "100000";
        when "1000010010010" => rgb <= "100000";
        when "1000010010011" => rgb <= "100000";
        when "1000010010100" => rgb <= "000000";
        when "1000010010111" => rgb <= "000000";
        when "1000010011000" => rgb <= "101000";
        when "1000010011001" => rgb <= "101000";
        when "1000010011010" => rgb <= "101000";
        when "1000010011011" => rgb <= "000000";
        when "1000010011110" => rgb <= "000000";
        when "1000010011111" => rgb <= "001010";
        when "1000010100000" => rgb <= "001010";
        when "1000010100001" => rgb <= "001010";
        when "1000010100010" => rgb <= "000000";
        when "1000010100011" => rgb <= "001010";
        when "1000010100100" => rgb <= "001010";
        when "1000010100101" => rgb <= "001010";
        when "1000010100110" => rgb <= "000000";
        when "1000010100111" => rgb <= "001010";
        when "1000010101000" => rgb <= "001010";
        when "1000010101001" => rgb <= "001010";
        when "1000010101010" => rgb <= "001010";
        when "1000010101011" => rgb <= "000000";
        when "1000010101100" => rgb <= "001010";
        when "1000010101101" => rgb <= "000000";
        when "1000010101110" => rgb <= "100110";
        when "1000010101111" => rgb <= "100110";
        when "1000010110000" => rgb <= "100110";
        when "1000010110001" => rgb <= "000000";
        when "1000010110100" => rgb <= "000000";
        when "1000010110101" => rgb <= "100110";
        when "1000010110110" => rgb <= "100110";
        when "1000010110111" => rgb <= "100110";
        when "1000010111000" => rgb <= "100110";
        when "1000010111001" => rgb <= "000000";
        when "1000010111100" => rgb <= "000000";
        when "1000010111101" => rgb <= "101000";
        when "1000010111110" => rgb <= "101000";
        when "1000010111111" => rgb <= "101000";
        when "1000011000000" => rgb <= "000000";
        when "1000100000110" => rgb <= "000000";
        when "1000100000111" => rgb <= "100000";
        when "1000100001000" => rgb <= "100000";
        when "1000100001001" => rgb <= "100000";
        when "1000100001010" => rgb <= "100000";
        when "1000100001011" => rgb <= "000000";
        when "1000100001100" => rgb <= "000000";
        when "1000100001101" => rgb <= "000000";
        when "1000100001110" => rgb <= "100000";
        when "1000100001111" => rgb <= "100000";
        when "1000100010000" => rgb <= "100000";
        when "1000100010001" => rgb <= "100000";
        when "1000100010010" => rgb <= "100000";
        when "1000100010011" => rgb <= "100000";
        when "1000100010100" => rgb <= "000000";
        when "1000100010111" => rgb <= "000000";
        when "1000100011000" => rgb <= "101000";
        when "1000100011001" => rgb <= "101000";
        when "1000100011010" => rgb <= "101000";
        when "1000100011011" => rgb <= "000000";
        when "1000100011110" => rgb <= "000000";
        when "1000100011111" => rgb <= "001010";
        when "1000100100000" => rgb <= "001010";
        when "1000100100001" => rgb <= "000000";
        when "1000100100010" => rgb <= "000000";
        when "1000100100011" => rgb <= "000000";
        when "1000100100100" => rgb <= "001010";
        when "1000100100101" => rgb <= "000000";
        when "1000100100110" => rgb <= "000000";
        when "1000100100111" => rgb <= "000000";
        when "1000100101000" => rgb <= "001010";
        when "1000100101001" => rgb <= "001010";
        when "1000100101010" => rgb <= "000000";
        when "1000100101011" => rgb <= "000000";
        when "1000100101100" => rgb <= "001010";
        when "1000100101101" => rgb <= "000000";
        when "1000100101110" => rgb <= "100110";
        when "1000100101111" => rgb <= "100110";
        when "1000100110000" => rgb <= "100110";
        when "1000100110001" => rgb <= "000000";
        when "1000100110100" => rgb <= "000000";
        when "1000100110101" => rgb <= "100110";
        when "1000100110110" => rgb <= "100110";
        when "1000100110111" => rgb <= "100110";
        when "1000100111000" => rgb <= "100110";
        when "1000100111001" => rgb <= "000000";
        when "1000100111100" => rgb <= "000000";
        when "1000100111101" => rgb <= "101000";
        when "1000100111110" => rgb <= "101000";
        when "1000100111111" => rgb <= "101000";
        when "1000101000000" => rgb <= "000000";
        when "1000110000101" => rgb <= "000000";
        when "1000110000110" => rgb <= "100000";
        when "1000110000111" => rgb <= "100000";
        when "1000110001000" => rgb <= "100000";
        when "1000110001001" => rgb <= "100000";
        when "1000110001010" => rgb <= "100000";
        when "1000110001011" => rgb <= "100000";
        when "1000110001100" => rgb <= "100000";
        when "1000110001101" => rgb <= "100000";
        when "1000110001110" => rgb <= "100000";
        when "1000110001111" => rgb <= "100000";
        when "1000110010000" => rgb <= "100000";
        when "1000110010001" => rgb <= "100000";
        when "1000110010010" => rgb <= "100000";
        when "1000110010011" => rgb <= "100000";
        when "1000110010100" => rgb <= "000000";
        when "1000110010111" => rgb <= "000000";
        when "1000110011000" => rgb <= "101000";
        when "1000110011001" => rgb <= "101000";
        when "1000110011010" => rgb <= "000000";
        when "1000110011110" => rgb <= "000000";
        when "1000110011111" => rgb <= "001010";
        when "1000110100000" => rgb <= "000000";
        when "1000110100001" => rgb <= "000000";
        when "1000110100011" => rgb <= "000000";
        when "1000110100100" => rgb <= "001010";
        when "1000110100101" => rgb <= "000000";
        when "1000110101000" => rgb <= "000000";
        when "1000110101001" => rgb <= "001010";
        when "1000110101010" => rgb <= "000000";
        when "1000110101100" => rgb <= "000000";
        when "1000110101101" => rgb <= "000000";
        when "1000110101110" => rgb <= "100110";
        when "1000110101111" => rgb <= "100110";
        when "1000110110000" => rgb <= "100110";
        when "1000110110001" => rgb <= "000000";
        when "1000110110101" => rgb <= "000000";
        when "1000110110110" => rgb <= "100110";
        when "1000110110111" => rgb <= "100110";
        when "1000110111000" => rgb <= "100110";
        when "1000110111001" => rgb <= "100110";
        when "1000110111010" => rgb <= "000000";
        when "1000110111100" => rgb <= "000000";
        when "1000110111101" => rgb <= "000000";
        when "1000110111110" => rgb <= "101000";
        when "1000110111111" => rgb <= "101000";
        when "1000111000000" => rgb <= "000000";
        when "1001000000110" => rgb <= "000000";
        when "1001000000111" => rgb <= "100000";
        when "1001000001000" => rgb <= "100000";
        when "1001000001001" => rgb <= "100000";
        when "1001000001010" => rgb <= "100000";
        when "1001000001011" => rgb <= "100000";
        when "1001000001100" => rgb <= "100000";
        when "1001000001101" => rgb <= "100000";
        when "1001000001110" => rgb <= "100000";
        when "1001000001111" => rgb <= "100000";
        when "1001000010000" => rgb <= "100000";
        when "1001000010001" => rgb <= "100000";
        when "1001000010010" => rgb <= "100000";
        when "1001000010011" => rgb <= "000000";
        when "1001000011000" => rgb <= "000000";
        when "1001000011001" => rgb <= "000000";
        when "1001000011111" => rgb <= "000000";
        when "1001000100000" => rgb <= "000000";
        when "1001000100100" => rgb <= "000000";
        when "1001000100101" => rgb <= "000000";
        when "1001000101001" => rgb <= "000000";
        when "1001000101101" => rgb <= "000000";
        when "1001000101110" => rgb <= "000000";
        when "1001000101111" => rgb <= "100110";
        when "1001000110000" => rgb <= "100110";
        when "1001000110001" => rgb <= "000000";
        when "1001000110101" => rgb <= "000000";
        when "1001000110110" => rgb <= "000000";
        when "1001000110111" => rgb <= "100110";
        when "1001000111000" => rgb <= "100110";
        when "1001000111001" => rgb <= "000000";
        when "1001000111010" => rgb <= "000000";
        when "1001000111101" => rgb <= "000000";
        when "1001000111110" => rgb <= "000000";
        when "1001000111111" => rgb <= "000000";
        when "1001010000110" => rgb <= "000000";
        when "1001010000111" => rgb <= "000000";
        when "1001010001000" => rgb <= "100000";
        when "1001010001001" => rgb <= "100000";
        when "1001010001010" => rgb <= "100000";
        when "1001010001011" => rgb <= "100000";
        when "1001010001100" => rgb <= "100000";
        when "1001010001101" => rgb <= "100000";
        when "1001010001110" => rgb <= "100000";
        when "1001010001111" => rgb <= "100000";
        when "1001010010000" => rgb <= "100000";
        when "1001010010001" => rgb <= "100000";
        when "1001010010010" => rgb <= "000000";
        when "1001010010011" => rgb <= "000000";
        when "1001010101110" => rgb <= "000000";
        when "1001010101111" => rgb <= "000000";
        when "1001010110000" => rgb <= "000000";
        when "1001010110001" => rgb <= "000000";
        when "1001010110111" => rgb <= "000000";
        when "1001010111000" => rgb <= "000000";
        when "1001100001000" => rgb <= "000000";
        when "1001100001001" => rgb <= "000000";
        when "1001100001010" => rgb <= "000000";
        when "1001100001011" => rgb <= "100000";
        when "1001100001100" => rgb <= "100000";
        when "1001100001101" => rgb <= "100000";
        when "1001100001110" => rgb <= "000000";
        when "1001100001111" => rgb <= "000000";
        when "1001100010000" => rgb <= "000000";
        when "1001100010001" => rgb <= "000000";
        when "1001110001011" => rgb <= "000000";
        when "1001110001100" => rgb <= "000000";
        when "1001110001101" => rgb <= "000000";
        when others => rgb <= "001000";
            end case;
   end process;
   position <= y_coord & x_coord;
end Behavioral;